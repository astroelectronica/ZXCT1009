.title KiCad schematic
.include "C:/AE/ZXCT1009/_models/BZX84C5V1.spice.txt"
.include "C:/AE/ZXCT1009/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/ZXCT1009/_models/CGJ4C2C0G2A101J060AA_p.mod"
.include "C:/AE/ZXCT1009/_models/FMMT597.spice.txt"
.include "C:/AE/ZXCT1009/_models/SMAZ15.spice.txt"
.include "C:/AE/ZXCT1009/_models/ZXCT1009.spice.txt"
R6 /PWR_OUT /SN {RLIM}
R5 /SN 0 {RTRAN}
I1 /PWR_OUT 0 PULSE( 0 {ILOAD} {TDELAY} {TR} {TF} {DUTY} {CYCLE} ) 
XU5 /PWR_IN /SN CGJ4C2C0G2A101J060AA_p
XU4 /SN /PWR_IN /COCM ZXCT1009F
R8 /PWR_IN /PWR_OUT {RSENSE2}
R7 /PWR_IN /PWR_OUT {RSENSE1}
R1 /OUT /FILTER {RFILTER}
XU2 /OUT 0 C2012C0G2A102J060AA_p
XU1 0 /OUT DI_BZX84C5V1
Q1 /FILTER /BASE /COCM FMMT597
R2 /FILTER 0 {RSET1}
R4 /FILTER 0 {RSET2}
R3 /BASE 0 {RBASE}
XU3 /BASE /PWR_IN SMAZ15
V1 /PWR_IN 0 {VSOURCE}
.end
